`timescale 1ns/1ns

`ifdef UVM_SIM
import uvm_pkg::*;
`include "uvm_macros.svh"
`endif

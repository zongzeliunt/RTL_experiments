`timescale 1ns/1ps

`ifdef UVM_SIM
import uvm_pkg::*;
`include "uvm_macros.svh"
`endif

`define LENGTH 4

interface Bus_if (input bit clk);
    wire reset;
    reg [3:0] data;
endinterface

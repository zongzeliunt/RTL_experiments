
	input [DATA_BITS - 1 : 0] input_data,
	output [DATA_BITS - 1 : 0] output_data,
	
	input wire read,
	input wire write,
	output wire empty,
	output wire full

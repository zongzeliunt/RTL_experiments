`timescale 1ns/1ns
import uvm_pkg::*;
`include "uvm_macros.svh"

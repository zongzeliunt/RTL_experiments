`timescale 1ns/1ps

`ifdef UVM_TB_SIM
import uvm_pkg::*;
`include "uvm_macros.svh"
`endif
